module cell (
  input x,
  output y
);

begin
endmodule
