module neuron (
  input [7:0]  D0, D1, D2, D3, D4, D5, D6, D7;
  output [7:0] Q;
);

   begin
      // empty module
endmodule // neuron


   
